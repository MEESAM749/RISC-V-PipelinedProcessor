module RISC_V_Processor ();

endmodule
